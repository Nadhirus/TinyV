module top;
  // Clock and reset signals
  logic clk;
  logic reset;


endmodule
